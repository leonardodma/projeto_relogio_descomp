library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 8;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  	constant NOP  : std_logic_vector(3 downto 0) := "0000";
	constant LDA  : std_logic_vector(3 downto 0) := "0001";
	constant SOMA : std_logic_vector(3 downto 0) := "0010";
	constant SUB  : std_logic_vector(3 downto 0) := "0011";
	constant LDI  : std_logic_vector(3 downto 0) := "0100";
	constant STA  : std_logic_vector(3 downto 0) := "0101";
	constant JMP  : std_logic_vector(3 downto 0) := "0110";
	constant JEQ  : std_logic_vector(3 downto 0) := "0111";
	constant CEQ  : std_logic_vector(3 downto 0) := "1000";
	constant JSR  : std_logic_vector(3 downto 0) := "1001";
	constant RET  : std_logic_vector(3 downto 0) := "1010";
  
  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  
tmp(0) := "0100000000000";	-- LDI $0				#Carrega o acumulador com o valor 0
tmp(1) := "0101100100000";	-- STA @288			#Armazena o valor do acumulador em HEX0
tmp(2) := "0101100100001";	-- STA @289			#Armazena o valor do acumulador em HEX1
tmp(3) := "0101100100010";	-- STA @290			#Armazena o valor do acumulador em HEX2
tmp(4) := "0101100100011";	-- STA @291			#Armazena o valor do acumulador em HEX3
tmp(5) := "0101100100100";	-- STA @292			#Armazena o valor do acumulador em HEX4
tmp(6) := "0101100100101";	-- STA @293			#Armazena o valor do acumulador em HEX5
tmp(7) := "0101100000000";	-- STA @256	    	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(8) := "0101100000001";	-- STA @257	    	#Armazena o valor do bit0 do acumulador no LDR8
tmp(9) := "0101100000010";	-- STA @258	    	#Armazena o valor do bit0 do acumulador no LDR9
tmp(10) := "0100000000000";	-- LDI $0				#Carrega o acumulador com o valor 0
tmp(11) := "0101000000000";	-- STA @0				#Armazena o valor do acumulador em MEM[0] (unidades)
tmp(12) := "0101000000001";	-- STA @1				#Armazena o valor do acumulador em MEM[1] (dezenas)
tmp(13) := "0101000000010";	-- STA @2				#Armazena o valor do acumulador em MEM[2] (centenas)
tmp(14) := "0100000000111";	-- LDI $7          	#Carrega o acumulador com o valor 7
tmp(15) := "0101000000011";	-- STA @3          	#Armazena o valor do acumulador em MEM[3] (LIMITE_UNID)
tmp(16) := "0101000000100";	-- STA @4          	#Armazena o valor do acumulador em MEM[4] (LIMITE_DEZ)
tmp(17) := "0101000000101";	-- STA @5          	#Armazena o valor do acumulador em MEM[5] (LIMITE_CENT)
tmp(18) := "0100000000000";	-- LDI $0          	#Carrega o acumulador com o valor 0
tmp(19) := "0101000000110";	-- STA @6          	#Armazena 0 ao acumulador em MEM[6] para comparacoes
tmp(20) := "0100000000001";	-- LDI $1          	#Carrega o acumulador com o valor 1
tmp(21) := "0101000000111";	-- STA @7          	#Armazena 1 ao acumulador em MEM[7] para incremento
tmp(22) := "0100000001010";	-- LDI $10         	#Carrega o acumulador com o valor 10
tmp(23) := "0101000001000";	-- STA @8          	#Armazena 10 ao acumulador em MEM[8] para comparacoes displays HEXs 
tmp(24) := "0100000000000";	-- LDI $0          	#Carrega o acumulador com o valor 0
tmp(25) := "0101000001001";	-- STA @9          	#Armazena 10 ao acumulador em MEM[9] para prosseguir ou não a contagem
tmp(26) := "0001101100000";	-- LDA @352
tmp(27) := "1000000001001";	-- CEQ @9
tmp(28) := "0111000011010";	-- JEQ FUNC_VERIFICA_KEY0
tmp(29) := "1001000100101";	-- JSR FUNC_INC_UNID
tmp(30) := "0001000000000";	-- LDA @0                
tmp(31) := "0101100100000";	-- STA @288                  
tmp(32) := "0001000000001";	-- LDA @1                
tmp(33) := "0101100100001";	-- STA @289 
tmp(34) := "0001000000010";	-- LDA @2                
tmp(35) := "0101100100010";	-- STA @290 
tmp(36) := "0110000011010";	-- JMP FUNC_VERIFICA_KEY0
tmp(37) := "0001000000000";	-- LDA @0    	#Armazena o valor MEM[0] no acumulador     
tmp(38) := "0010000000111";	-- SOMA @7                  	#Soma o valor do acumulador com o MEM[7]                 
tmp(39) := "1000000001000";	-- CEQ @8		             	#Compara o valor do acumulador com o MEM[8]
tmp(40) := "0111000101011";	-- JEQ FUNC_INC_DEZENA      	#Se for 0 incrementa DEZENA, se não incrementa UNID
tmp(41) := "0101000000000";	-- STA @0
tmp(42) := "1010000000000";	-- RET
tmp(43) := "0001000000001";	-- LDA @1  	#Armazena o valor MEM[1] no acumulador 
tmp(44) := "0010000000111";	-- SOMA @7                  	#Soma o valor do acumulador com o MEM[7]                 
tmp(45) := "1000000001000";	-- CEQ @8		             	#Compara o valor do acumulador com o MEM[8]
tmp(46) := "0111000110001";	-- JEQ FUNC_INC_CENTENA      	#Se for 0 incrementa CENTENA, se não incrementa DEZENA
tmp(47) := "0101000000001";	-- STA @1
tmp(48) := "1010000000000";	-- RET
tmp(49) := "0001000000010";	-- LDA @2  	#Armazena o valor MEM[2] no acumulador 
tmp(50) := "0010000000111";	-- SOMA @7                   	#Soma o valor do acumulador com o MEM[7]                 
tmp(51) := "1000000001000";	-- CEQ @8		              	#Compara o valor do acumulador com o MEM[8]
tmp(52) := "0111000000000";	-- JEQ FUNC_SETUP            	#Se for 0 incrementa CENTENA, se não incrementa CENTENA
tmp(53) := "0101000000010";	-- STA @2
tmp(54) := "1010000000000";	-- RET


        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;